`ifndef CONFIG
`define CONFIG

`define DATA_WIDTH 32
`define INST_WIDTH 32


`endif 